//Copyright (C)2014-2021 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//GOWIN Version: V1.9.8
//Part Number: GW1N-LV9QN88C6/I5
//Device: GW1N-9
//Created Time: Fri Nov 12 14:09:56 2021

module bootram_2kx8_1 (dout, clk, oce, ce, reset, wre, ad, din);

output [7:0] dout;
input clk;
input oce;
input ce;
input reset;
input wre;
input [10:0] ad;
input [7:0] din;

wire [23:0] sp_inst_0_dout_w;
wire gw_gnd;

assign gw_gnd = 1'b0;

SP sp_inst_0 (
    .DO({sp_inst_0_dout_w[23:0],dout[7:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,gw_gnd}),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[7:0]})
);

defparam sp_inst_0.READ_MODE = 1'b0;
defparam sp_inst_0.WRITE_MODE = 2'b00;
defparam sp_inst_0.BIT_WIDTH = 8;
defparam sp_inst_0.BLK_SEL = 3'b000;
defparam sp_inst_0.RESET_MODE = "SYNC";
defparam sp_inst_0.INIT_RAM_00 = 256'h252523232220000120222426282A2C2E20222426282A2C2E0000000000000000;
defparam sp_inst_0.INIT_RAM_01 = 256'h2005260E8515010515F00520088515051581811100012F2F2E2E282827272626;
defparam sp_inst_0.INIT_RAM_02 = 256'h0747A6A817A0A40707A207072E20222426282A2C2E2022242601000001F02580;
defparam sp_inst_0.INIT_RAM_03 = 256'h58A6A886A64C0747A6A820060758A6A886A64C0747A6A820060758A6A886A64C;
defparam sp_inst_0.INIT_RAM_04 = 256'h47A6A820060758A6A886A64C0747A6A820060758A6A886A64C0747A6A8200607;
defparam sp_inst_0.INIT_RAM_05 = 256'hA6A886A64C0747A6A820060758A6A886A64C0747A6A820060758A6A886A64C07;
defparam sp_inst_0.INIT_RAM_06 = 256'h07A007A0070758A6A886A64C0747A6A820060758A6A886A64C0747A6A8200758;
defparam sp_inst_0.INIT_RAM_07 = 256'h070717A007079847A08A07060605070717A007079847A08C07060605070717A0;
defparam sp_inst_0.INIT_RAM_08 = 256'h07060605070717A007079847A08607060605070717A007079847A08807060605;
defparam sp_inst_0.INIT_RAM_09 = 256'h1A17248717A007A007079847A08407060605070717A007A007A007079847A082;
defparam sp_inst_0.INIT_RAM_0A = 256'h8E0686072020200F030F09020A0C04040B060B080709268D808E8A19871D101E;
defparam sp_inst_0.INIT_RAM_0B = 256'h0820458676D68620458676D60420458676D68220458676D6004586D627984720;
defparam sp_inst_0.INIT_RAM_0C = 256'h2727279847208006070620052020208E20C787F70C20468676D68A20458676D6;
defparam sp_inst_0.INIT_RAM_0D = 256'h47A0A0F09047A0A0F09E47A0A0F09C47A0A080A78797E087202020E4F776868C;
defparam sp_inst_0.INIT_RAM_0E = 256'hD6479605058708B72E23F020C727F020C727F020C727F020C727F020C727F092;
defparam sp_inst_0.INIT_RAM_0F = 256'h200685852006252818081AC70526108C0685000D0D0ACD06050C908580C796C7;
defparam sp_inst_0.INIT_RAM_10 = 256'hD68020458676D60E20488676D68C20458676D60A20488676D6884586D60318C6;
defparam sp_inst_0.INIT_RAM_11 = 256'h804586560E18C6200E8506202025202006204686F38420458676D60220488676;
defparam sp_inst_0.INIT_RAM_12 = 256'h76560A2045867656882045867656062045867656842045867656022045867656;
defparam sp_inst_0.INIT_RAM_13 = 256'h76D68C20458676D60A4586D618C62008850620202520200E2046867E8C204586;
defparam sp_inst_0.INIT_RAM_14 = 256'h20C787F70620468676D68420458676D60220458676D68020458676D60E204586;
defparam sp_inst_0.INIT_RAM_15 = 256'h76D6922020458676D6144586D6279A472020F098472020F020C727F020202088;
defparam sp_inst_0.INIT_RAM_16 = 256'h2020468676D69A2020458676D61C2020458676D69E2020458676D61020204586;
defparam sp_inst_0.INIT_RAM_17 = 256'h982020458676D61A2020488676D69C4586D60312C62020F020962020C787F718;
defparam sp_inst_0.INIT_RAM_18 = 256'h204686F3902020458676D6122020488676D6942020458676D6162020488676D6;
defparam sp_inst_0.INIT_RAM_19 = 256'h2020458676D6162020458676D6982020458676D61A4586D610C62020F0201E20;
defparam sp_inst_0.INIT_RAM_1A = 256'h2020F0209C2020C787F71E2020468676D6902020458676D6122020458676D694;
defparam sp_inst_0.INIT_RAM_1B = 256'h458676561E2020458676569020204586765612202045867656944586560E1AC6;
defparam sp_inst_0.INIT_RAM_1C = 256'h9447A0A0F08E85F02016202046867E982020458676561A2020458676569C2020;
defparam sp_inst_0.INIT_RAM_1D = 256'h5F20205F2020205F20786D6878736E7873790A07070707070780F09647A0A0F0;
defparam sp_inst_0.INIT_RAM_1E = 256'h207C005F20205F297C7C5F7C0A5C2F5F205F7C297C0A5F20205F5F5F29207C00;
defparam sp_inst_0.INIT_RAM_1F = 256'h000000000064393531006E6F20614F0A6F205468202020200A5F2F5C5F5F5F7C;
defparam sp_inst_0.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

endmodule //bootram_2kx8_1
