//Copyright (C)2014-2021 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//GOWIN Version: V1.9.8
//Part Number: GW1N-LV9QN88C6/I5
//Device: GW1N-9
//Created Time: Wed Nov 10 21:40:34 2021

module bootram_4k (dout, clk, oce, ce, reset, wre, ad, din);

output [31:0] dout;
input clk;
input oce;
input ce;
input reset;
input wre;
input [9:0] ad;
input [31:0] din;

wire [15:0] sp_inst_0_dout_w;
wire [15:0] sp_inst_1_dout_w;
wire gw_vcc;
wire gw_gnd;

assign gw_vcc = 1'b1;
assign gw_gnd = 1'b0;

SP sp_inst_0 (
    .DO({sp_inst_0_dout_w[15:0],dout[15:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,gw_gnd}),
    .AD({ad[9:0],gw_gnd,gw_gnd,gw_vcc,gw_vcc}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]})
);

defparam sp_inst_0.READ_MODE = 1'b0;
defparam sp_inst_0.WRITE_MODE = 2'b00;
defparam sp_inst_0.BIT_WIDTH = 16;
defparam sp_inst_0.BLK_SEL = 3'b000;
defparam sp_inst_0.RESET_MODE = "SYNC";
defparam sp_inst_0.INIT_RAM_00 = 256'h202322232423262328232A232C232E230013001300130013001300130013006F;
defparam sp_inst_0.INIT_RAM_01 = 256'h25832503238323032283208300EF0113202322232423262328232A232C232E23;
defparam sp_inst_0.INIT_RAM_02 = 256'h0513011381931197007301132F832F032E832E03288328032783270326832603;
defparam sp_inst_0.INIT_RAM_03 = 256'h0113F06F250380E72023051326830E63059301130513F06F0513202308630593;
defparam sp_inst_0.INIT_RAM_04 = 256'h07930737A0230713A0230713A0230713A22307132423262307B70113006F00EF;
defparam sp_inst_0.INIT_RAM_05 = 256'h0593079307130737A023071307B798E34783A02380630713061306B705930713;
defparam sp_inst_0.INIT_RAM_06 = 256'h061306B70593071307930737A023071307B798E34783A0238E630713061306B7;
defparam sp_inst_0.INIT_RAM_07 = 256'h8A630713061306B70593079307130737A023071307B798E34783A0238C630713;
defparam sp_inst_0.INIT_RAM_08 = 256'h4783A0238E630713061306B70593071307930737A023071307B798E34783A023;
defparam sp_inst_0.INIT_RAM_09 = 256'h80630713061306B70593079307130737A0230713A0230713A023071307B798E3;
defparam sp_inst_0.INIT_RAM_0A = 256'h041306930E1305938F938093A0230FB7071300B7A023071307B798E34783A023;
defparam sp_inst_0.INIT_RAM_0B = 256'h0E63061307138613A023A023A023A023A0230F37051308130893029303130393;
defparam sp_inst_0.INIT_RAM_0C = 256'h0CE3A7032773277318E34703A0230263061386130713A0230E9318E34703A023;
defparam sp_inst_0.INIT_RAM_0D = 256'h4783A023A023F06F92E38E9304630E630863A023A023A023E463771376130613;
defparam sp_inst_0.INIT_RAM_0E = 256'h9EE34783A023A023F06F9CE34783A023A023F06F9AE34783A023A023F06F98E3;
defparam sp_inst_0.INIT_RAM_0F = 256'h2703F06F202347132703F06F1AE34703A023A023F06F16E34703A023A023F06F;
defparam sp_inst_0.INIT_RAM_10 = 256'h9AE34783A023A023F06F98E34783A023A023F06F202347132703F06F20234713;
defparam sp_inst_0.INIT_RAM_11 = 256'h5F5F295F205F7C20000A5F5F202020205F5F20202020205F5F5F20208067F06F;
defparam sp_inst_0.INIT_RAM_12 = 256'h7C200A7C5C202F205F5F205F5F5F7C20295F7C200A7C5F20205F20205F5F5F5F;
defparam sp_inst_0.INIT_RAM_13 = 256'h5C205F5F5F5F5F5F7C5F20207C20000A5F7C2029207C5F5F295F7C5F7C205F5F;
defparam sp_inst_0.INIT_RAM_14 = 256'h6F433A65745350530A4B6F6E206754206863206E2020202020200A7C5F5F2F5F;
defparam sp_inst_0.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000206E61;
defparam sp_inst_0.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_1 (
    .DO({sp_inst_1_dout_w[15:0],dout[31:16]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,gw_gnd}),
    .AD({ad[9:0],gw_gnd,gw_gnd,gw_vcc,gw_vcc}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[31:16]})
);

defparam sp_inst_1.READ_MODE = 1'b0;
defparam sp_inst_1.WRITE_MODE = 2'b00;
defparam sp_inst_1.BIT_WIDTH = 16;
defparam sp_inst_1.BLK_SEL = 3'b000;
defparam sp_inst_1.RESET_MODE = "SYNC";
defparam sp_inst_1.INIT_RAM_00 = 256'hFED1FEC1FEB1FEA1FE71FE61FE51FE1100000000000000000000000000000B00;
defparam sp_inst_1.INIT_RAM_01 = 256'h028102C103010341038103C13E00FC01FDF1FDE1FDD1FDC1FD11FD01FCF1FCE1;
defparam sp_inst_1.INIT_RAM_02 = 256'h54807500C98100003020040100010041008100C101010141018101C102010241;
defparam sp_inst_1.INIT_RAM_03 = 256'h0041FE5F0001000600A10045000500B55480FFC15480FF5F0045000500B55480;
defparam sp_inst_1.INIT_RAM_04 = 256'h0200000000E7020000E700A000E700D000E7002000810011C000FF0100000080;
defparam sp_inst_1.INIT_RAM_05 = 256'h00A007C04717000000E70200C000FE07000700F622B7001700D0C00000A04497;
defparam sp_inst_1.INIT_RAM_06 = 256'h00D0C00000A0499707C0000000E70200C000FE07000700F61EB7001700D0C000;
defparam sp_inst_1.INIT_RAM_07 = 256'h1AB7001700D0C00000A007C04BD7000000E70200C000FE07000700F61CB70017;
defparam sp_inst_1.INIT_RAM_08 = 256'h000700F61EB7001700D0C00000A04E5707C0000000E70200C000FE07000700F6;
defparam sp_inst_1.INIT_RAM_09 = 256'h1AB7001700D0C00000A0020050D7000000E7020000E700A000E700D0C000FE07;
defparam sp_inst_1.INIT_RAM_0A = 256'h053000A000D000D053DF531000E7000000A0000000E700D0C000FE07000700F6;
defparam sp_inst_1.INIT_RAM_0B = 256'h0CD7001605000000008700D701C700D701C7800003700390038005D0FFF00430;
defparam sp_inst_1.INIT_RAM_0C = 256'hFE670007C000C000FE07000600E70AD70016000F06F0007700A0FE07000600E7;
defparam sp_inst_1.INIT_RAM_0D = 256'h000700F600C6F6DFFA0EFFFE08A709070B1700D700B700E700C20FF70FF6FDF7;
defparam sp_inst_1.INIT_RAM_0E = 256'hE207000700F600C6E29FE007000700F600C6E05FDE07000700F600C6DE1FDC07;
defparam sp_inst_1.INIT_RAM_0F = 256'h000FEE5F00EF0017000FF25FF007000600E700B7F5DFF407000600E700B7E4DF;
defparam sp_inst_1.INIT_RAM_10 = 256'hDE07000700F600C6E61FE407000700F600C6EC5F00EF0027000FED5F00EF0047;
defparam sp_inst_1.INIT_RAM_11 = 256'h5F205F20285C202000005F5F20202020205F5F202020202020205F5F0000E05F;
defparam sp_inst_1.INIT_RAM_12 = 256'h20200000207C5F205C205F5C202F202F7C207C2000005F5F2F205F5F7C5F202F;
defparam sp_inst_1.INIT_RAM_13 = 256'h5F5F2F5F5F2F5F5C5F5C7C207C5F00005F5F207C5F2820297C20282028207C2F;
defparam sp_inst_1.INIT_RAM_14 = 256'h6D6D000A746120490000392D614E6E616565694C4F202020202000005F5F5C20;
defparam sp_inst_1.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000003E64;
defparam sp_inst_1.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

endmodule //bootram_4k
