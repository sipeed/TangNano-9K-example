//Copyright (C)2014-2021 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//GOWIN Version: V1.9.8
//Part Number: GW1N-LV9QN88C6/I5
//Device: GW1N-9
//Created Time: Fri Nov 12 14:10:06 2021

module bootram_2kx8_2 (dout, clk, oce, ce, reset, wre, ad, din);

output [7:0] dout;
input clk;
input oce;
input ce;
input reset;
input wre;
input [10:0] ad;
input [7:0] din;

wire [23:0] sp_inst_0_dout_w;
wire gw_gnd;

assign gw_gnd = 1'b0;

SP sp_inst_0 (
    .DO({sp_inst_0_dout_w[23:0],dout[7:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,gw_gnd}),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[7:0]})
);

defparam sp_inst_0.READ_MODE = 1'b0;
defparam sp_inst_0.WRITE_MODE = 2'b00;
defparam sp_inst_0.BIT_WIDTH = 8;
defparam sp_inst_0.BLK_SEL = 3'b000;
defparam sp_inst_0.RESET_MODE = "SYNC";
defparam sp_inst_0.INIT_RAM_00 = 256'h81C1014181C15001F1E1D1C11101F1E1D1C1B1A1716151110000000000000000;
defparam sp_inst_0.INIT_RAM_01 = 256'hA14505B58500C145005F4505B5050045000101002001014181C1014181C10141;
defparam sp_inst_0.INIT_RAM_02 = 256'hF70F070700E7E7F000E79000B1A19181716151413121918111010080411F0106;
defparam sp_inst_0.INIT_RAM_03 = 256'hD707D71607D7F70F0707D7D000D707D71607D7F70F0707D7E000D707D71607D7;
defparam sp_inst_0.INIT_RAM_04 = 256'h0F0707D7F000D707D71607D7F70F0707D77000D707D71607D7F70F0707D7B000;
defparam sp_inst_0.INIT_RAM_05 = 256'h07D71607D7F70F0707D7F000D707D71607D7F70F0707D7F000D707D71607D7F7;
defparam sp_inst_0.INIT_RAM_06 = 256'h00E7A0E7D000D707D71607D7F70F0707D7F000D707D71607D7F70F07070700D7;
defparam sp_inst_0.INIT_RAM_07 = 256'hC0D700E700000707F6B717D000A057C000E700000707F6B717D000A000D700E7;
defparam sp_inst_0.INIT_RAM_08 = 256'h17D000A0C09700E700000707F6B717D000A017C000E700000707F6B717D000A0;
defparam sp_inst_0.INIT_RAM_09 = 256'h0000F15700E7A0E7D0000707F6B717D000A0001700E700E7A0E7D0000707F6B7;
defparam sp_inst_0.INIT_RAM_0A = 256'hD7160AF0976777000160D0F030300090A0A0D0D00019F19DC0CE5A0017000000;
defparam sp_inst_0.INIT_RAM_0B = 256'hD5B706CEF6C7D5A706CEF607D5B706CEF647D5A706CEF687D506CEC7040706F7;
defparam sp_inst_0.INIT_RAM_0C = 256'h0700000706F7D716F00947A0D717F7D7C707FEF7D6B706CEF647D5A706CEF687;
defparam sp_inst_0.INIT_RAM_0D = 256'h07F6C61F0707F6C6DF0707F6C69F0707F6C60707F027FF07D717F7C9F7F6F757;
defparam sp_inst_0.INIT_RAM_0E = 256'h17F6D705011740B920001FF417041FF427041FF447041FF487041FF407045F07;
defparam sp_inst_0.INIT_RAM_0F = 256'hC7D6150D8790200008F865C74505E61C1615CDBD010D0C0000016515F5C757C7;
defparam sp_inst_0.INIT_RAM_10 = 256'h83D50706CEF6C3D8B706CEF603D50706CEF643D8B706CEF683D506CEC3780605;
defparam sp_inst_0.INIT_RAM_11 = 256'hD506CECEC50605C7D615E097D78117C7D6B7067EF3D50706CEF643D8B706CEF6;
defparam sp_inst_0.INIT_RAM_12 = 256'hF64ED5B706CEF68ED5A706CEF6CED5B706CEF60ED5A706CEF64ED5B706CEF68E;
defparam sp_inst_0.INIT_RAM_13 = 256'hF647D5A706CEF687D506CEC70605C7D6158087D7C117C7D6B706CEFED5A706CE;
defparam sp_inst_0.INIT_RAM_14 = 256'hC707FEF7D6B706CEF647D5A706CEF687D5B706CEF6C7D5A706CEF607D5B706CE;
defparam sp_inst_0.INIT_RAM_15 = 256'hF647D5A71706CEF687D506CEC7040706F7171F0706F7175FF407045FD717F7D7;
defparam sp_inst_0.INIT_RAM_16 = 256'hB71706CEF647D5A71706CEF687D5B71706CEF6C7D5A71706CEF607D5B71706CE;
defparam sp_inst_0.INIT_RAM_17 = 256'hD5071706CEF643D8B71706CEF683D506CEC3780605C7175F17D7C71707FEF7D6;
defparam sp_inst_0.INIT_RAM_18 = 256'h17067EF3D5071706CEF643D8B71706CEF683D5071706CEF6C3D8B71706CEF603;
defparam sp_inst_0.INIT_RAM_19 = 256'hA71706CEF607D5B71706CEF647D5A71706CEF687D506CEC70605C7175F17D6B7;
defparam sp_inst_0.INIT_RAM_1A = 256'hC7171F17D7C71707FEF7D6B71706CEF647D5A71706CEF687D5B71706CEF6C7D5;
defparam sp_inst_0.INIT_RAM_1B = 256'h06CEF6CED5B71706CEF60ED5A71706CEF64ED5B71706CEF68ED506CECEC50605;
defparam sp_inst_0.INIT_RAM_1C = 256'h0707F6C68F05F55F17D6B71706CEFED5A71706CEF64ED5B71706CEF68ED5A717;
defparam sp_inst_0.INIT_RAM_1D = 256'h5F20205F202020205F003A6B003A73003A630000000000000000CF0707F6C68F;
defparam sp_inst_0.INIT_RAM_1E = 256'h205F005F7C28292020202F20007C20205C2F2F2020005F205F5F2F20205C2000;
defparam sp_inst_0.INIT_RAM_1F = 256'h00000000006561363200646D007420002D4E61654C202020005F205F5F2F5C5C;
defparam sp_inst_0.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

endmodule //bootram_2kx8_2
