//Copyright (C)2014-2021 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//GOWIN Version: V1.9.8
//Part Number: GW1N-LV9QN88C6/I5
//Device: GW1N-9
//Created Time: Fri Nov 12 14:10:17 2021

module bootram_2kx8_3 (dout, clk, oce, ce, reset, wre, ad, din);

output [7:0] dout;
input clk;
input oce;
input ce;
input reset;
input wre;
input [10:0] ad;
input [7:0] din;

wire [23:0] sp_inst_0_dout_w;
wire gw_gnd;

assign gw_gnd = 1'b0;

SP sp_inst_0 (
    .DO({sp_inst_0_dout_w[23:0],dout[7:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,gw_gnd}),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[7:0]})
);

defparam sp_inst_0.READ_MODE = 1'b0;
defparam sp_inst_0.WRITE_MODE = 2'b00;
defparam sp_inst_0.BIT_WIDTH = 8;
defparam sp_inst_0.BLK_SEL = 3'b000;
defparam sp_inst_0.RESET_MODE = "SYNC";
defparam sp_inst_0.INIT_RAM_00 = 256'h02020303030363FCFDFDFDFDFDFDFCFCFEFEFEFEFEFEFEFE000000000000000B;
defparam sp_inst_0.INIT_RAM_01 = 256'h00000000F000FFF100FF000000F300F300C17400300400000000010101010202;
defparam sp_inst_0.INIT_RAM_02 = 256'h2300FFFE0000000380000EC011131313131313131315141414EB000000FE0000;
defparam sp_inst_0.INIT_RAM_03 = 256'hFEFFFE00FF002300FFFE000380FEFFFE00FF002300FFFE000380FEFFFE00FF00;
defparam sp_inst_0.INIT_RAM_04 = 256'h00FFFE000280FEFFFE00FF002300FFFE000380FEFFFE00FF002300FFFE000380;
defparam sp_inst_0.INIT_RAM_05 = 256'hFFFE00FF002300FFFE000380FEFFFE00FF002300FFFE000180FEFFFE00FF0023;
defparam sp_inst_0.INIT_RAM_06 = 256'h0200000000C0FEFFFE00FF002300FFFE000380FEFFFE00FF002300FFFE0080FE;
defparam sp_inst_0.INIT_RAM_07 = 256'h07F2000002C0FE00002E0000C000F007000002C0FE0000300000C00002ED0000;
defparam sp_inst_0.INIT_RAM_08 = 256'h0000C00007F7000002C0FE00002A0000C000F507000002C0FE00002C0000C000;
defparam sp_inst_0.INIT_RAM_09 = 256'h000000EC0000000000C0FE00001A0000C00002FA00000200000000C0FE000020;
defparam sp_inst_0.INIT_RAM_0A = 256'h5200000400010110110005FF0404800400000000C0FD00EBE9FDFC00ED000000;
defparam sp_inst_0.INIT_RAM_0B = 256'h5400000000005400000000015400000000015400000000015400000100FE0000;
defparam sp_inst_0.INIT_RAM_0C = 256'h00C0C0FE00004400060001000001005400000000540000000000540000000000;
defparam sp_inst_0.INIT_RAM_0D = 256'h000000D3D2000000D0CE000000CECC000000000000007CFD000100000F0FFDFE;
defparam sp_inst_0.INIT_RAM_0E = 256'h01000000010A0112C0C0E1000000E2000000E3000000E4000000E5000100D5D4;
defparam sp_inst_0.INIT_RAM_0F = 256'h003A00000107C0C0F8FFFE000000FF000000F000110000000001FE0000000000;
defparam sp_inst_0.INIT_RAM_10 = 256'h003C01000000003A00000000013A01000000013A00000000013A00000140FE00;
defparam sp_inst_0.INIT_RAM_11 = 256'h4A00000141FE000048000600000001003C000000003C01000000003C00000000;
defparam sp_inst_0.INIT_RAM_12 = 256'h00004A00000000004A00000000004A00000000014A00000000014A0000000001;
defparam sp_inst_0.INIT_RAM_13 = 256'h00012C00000000012C000001FE00002C000601000001004A000001004A000000;
defparam sp_inst_0.INIT_RAM_14 = 256'h000000002E00000000002E00000000002E00000000002E00000000012C000000;
defparam sp_inst_0.INIT_RAM_15 = 256'h0001AC000100000001AC00000100AA000001BCBA000001AC000200AD0001002E;
defparam sp_inst_0.INIT_RAM_16 = 256'h000100000000AA000100000000AA000100000000AA000100000001AC00010000;
defparam sp_inst_0.INIT_RAM_17 = 256'hC4010100000001C4000100000001C400000140C4000001AA01AA0001000000AA;
defparam sp_inst_0.INIT_RAM_18 = 256'h01000000C4010100000000C4000100000000C4010100000000C4000100000001;
defparam sp_inst_0.INIT_RAM_19 = 256'h000100000001D2000100000001D2000100000001D2000001D2000001C301C200;
defparam sp_inst_0.INIT_RAM_1A = 256'h0001D101D00001000000D0000100000000D2000100000000D2000100000000D2;
defparam sp_inst_0.INIT_RAM_1B = 256'h00000000B4000100000001B6000100000001B6000100000001B600000141B400;
defparam sp_inst_0.INIT_RAM_1C = 256'hE4000000FEEEFFB401B40001000100B4000100000000B4000100000000B40001;
defparam sp_inst_0.INIT_RAM_1D = 256'h5F2020205F2020205F00207300207400206C0000000000000000DFDE000000E5;
defparam sp_inst_0.INIT_RAM_1E = 256'h7C7C005F205F207C28287C2000205F5C5F20207C7C005F2F5F7C205F5F282000;
defparam sp_inst_0.INIT_RAM_1F = 256'h000000000066623733003E6D0065530039616E65694F2020005F5C5F2F5F5F5F;
defparam sp_inst_0.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

endmodule //bootram_2kx8_3
